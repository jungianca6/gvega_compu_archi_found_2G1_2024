module calculadoraFPGA (
		input logic a,b,c,d,
		output logic [2:0] resultado,
		output logic [3:0] display
);


	
endmodule